//==============================================================================
// Module name: silde
// Author     : momo
// E-mail     : 1345238761@qq.com
// Create date: 2019.7.8
// Description: idle for reset
// -------------------------------------------------
// Modification log here:
// Author     :
// Date       : 
// Message    :
//==============================================================================
module silde
(
  input               clk,
  input               rstn,

  input               en_idle
);

endmodule