module resetn
(
  input   SW1,
  output  rstn
);

  assign rstn = SW1;

endmodule