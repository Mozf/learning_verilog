//==============================================================================
// Module name: floor
// Author     : momo
// E-mail     : 1345238761@qq.com
// Create date: 2019.7.30
// Description: 
// -------------------------------------------------
// Modification log here:
// Author     :
// Date       : 
// Message    :
//==============================================================================
module floor
(
  input clk,
  input rstn,

  output reg  LED4_R,
  output reg  LED4_G,
  output reg  LED4_B,
);

endmodule